///////////////////////////////////////////////////////////////////////////////////////////////////////////////
//  Author : Sachin
//  Description :  
///////////////////////////////////////////////////////////////////////////////////////////////////////////////

module mux_2_1 (
        input wire in_0,
        input wire in_1,
        input wire sel,

        output logic out
);

assign out = sel ? in_1 : in_0;

endmodule
